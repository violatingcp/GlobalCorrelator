library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pf_constants is

  constant N_PF_IP_CORE_IN_CHANS : natural  := 112;
  constant N_PF_IP_CORE_OUT_CHANS : natural := 112;
  constant N_IN_CHANS  : natural := 112;
  constant N_OUT_CHANS : natural := 112;
  constant PAYLOAD_LATENCY : natural := 25;
  
end;
    
